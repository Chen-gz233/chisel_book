module RAM_1(
  input        clock,
  input        reset,
  input  [7:0] io_in_addr,
  input  [7:0] io_in_data,
  input        io_in_en,
  output [7:0] io_out_data,
  output       io_out_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] fifo_0; // @[main.scala 23:23]
  reg [7:0] fifo_1; // @[main.scala 23:23]
  reg [7:0] fifo_2; // @[main.scala 23:23]
  reg [7:0] fifo_3; // @[main.scala 23:23]
  reg [7:0] fifo_4; // @[main.scala 23:23]
  reg [7:0] fifo_5; // @[main.scala 23:23]
  reg [7:0] fifo_6; // @[main.scala 23:23]
  reg [7:0] fifo_7; // @[main.scala 23:23]
  reg [7:0] fifo_8; // @[main.scala 23:23]
  reg [7:0] fifo_9; // @[main.scala 23:23]
  reg [7:0] fifo_10; // @[main.scala 23:23]
  reg [7:0] fifo_11; // @[main.scala 23:23]
  reg [7:0] fifo_12; // @[main.scala 23:23]
  reg [7:0] fifo_13; // @[main.scala 23:23]
  reg [7:0] fifo_14; // @[main.scala 23:23]
  reg [7:0] fifo_15; // @[main.scala 23:23]
  reg [7:0] fifo_16; // @[main.scala 23:23]
  reg [7:0] fifo_17; // @[main.scala 23:23]
  reg [7:0] fifo_18; // @[main.scala 23:23]
  reg [7:0] fifo_19; // @[main.scala 23:23]
  reg [7:0] fifo_20; // @[main.scala 23:23]
  reg [7:0] fifo_21; // @[main.scala 23:23]
  reg [7:0] fifo_22; // @[main.scala 23:23]
  reg [7:0] fifo_23; // @[main.scala 23:23]
  reg [7:0] fifo_24; // @[main.scala 23:23]
  reg [7:0] fifo_25; // @[main.scala 23:23]
  reg [7:0] fifo_26; // @[main.scala 23:23]
  reg [7:0] fifo_27; // @[main.scala 23:23]
  reg [7:0] fifo_28; // @[main.scala 23:23]
  reg [7:0] fifo_29; // @[main.scala 23:23]
  reg [7:0] fifo_30; // @[main.scala 23:23]
  reg [7:0] fifo_31; // @[main.scala 23:23]
  reg [7:0] fifo_32; // @[main.scala 23:23]
  reg [7:0] fifo_33; // @[main.scala 23:23]
  reg [7:0] fifo_34; // @[main.scala 23:23]
  reg [7:0] fifo_35; // @[main.scala 23:23]
  reg [7:0] fifo_36; // @[main.scala 23:23]
  reg [7:0] fifo_37; // @[main.scala 23:23]
  reg [7:0] fifo_38; // @[main.scala 23:23]
  reg [7:0] fifo_39; // @[main.scala 23:23]
  reg [7:0] fifo_40; // @[main.scala 23:23]
  reg [7:0] fifo_41; // @[main.scala 23:23]
  reg [7:0] fifo_42; // @[main.scala 23:23]
  reg [7:0] fifo_43; // @[main.scala 23:23]
  reg [7:0] fifo_44; // @[main.scala 23:23]
  reg [7:0] fifo_45; // @[main.scala 23:23]
  reg [7:0] fifo_46; // @[main.scala 23:23]
  reg [7:0] fifo_47; // @[main.scala 23:23]
  reg [7:0] fifo_48; // @[main.scala 23:23]
  reg [7:0] fifo_49; // @[main.scala 23:23]
  reg [7:0] fifo_50; // @[main.scala 23:23]
  reg [7:0] fifo_51; // @[main.scala 23:23]
  reg [7:0] fifo_52; // @[main.scala 23:23]
  reg [7:0] fifo_53; // @[main.scala 23:23]
  reg [7:0] fifo_54; // @[main.scala 23:23]
  reg [7:0] fifo_55; // @[main.scala 23:23]
  reg [7:0] fifo_56; // @[main.scala 23:23]
  reg [7:0] fifo_57; // @[main.scala 23:23]
  reg [7:0] fifo_58; // @[main.scala 23:23]
  reg [7:0] fifo_59; // @[main.scala 23:23]
  reg [7:0] fifo_60; // @[main.scala 23:23]
  reg [7:0] fifo_61; // @[main.scala 23:23]
  reg [7:0] fifo_62; // @[main.scala 23:23]
  reg [7:0] fifo_63; // @[main.scala 23:23]
  reg [7:0] fifo_64; // @[main.scala 23:23]
  reg [7:0] fifo_65; // @[main.scala 23:23]
  reg [7:0] fifo_66; // @[main.scala 23:23]
  reg [7:0] fifo_67; // @[main.scala 23:23]
  reg [7:0] fifo_68; // @[main.scala 23:23]
  reg [7:0] fifo_69; // @[main.scala 23:23]
  reg [7:0] fifo_70; // @[main.scala 23:23]
  reg [7:0] fifo_71; // @[main.scala 23:23]
  reg [7:0] fifo_72; // @[main.scala 23:23]
  reg [7:0] fifo_73; // @[main.scala 23:23]
  reg [7:0] fifo_74; // @[main.scala 23:23]
  reg [7:0] fifo_75; // @[main.scala 23:23]
  reg [7:0] fifo_76; // @[main.scala 23:23]
  reg [7:0] fifo_77; // @[main.scala 23:23]
  reg [7:0] fifo_78; // @[main.scala 23:23]
  reg [7:0] fifo_79; // @[main.scala 23:23]
  reg [7:0] fifo_80; // @[main.scala 23:23]
  reg [7:0] fifo_81; // @[main.scala 23:23]
  reg [7:0] fifo_82; // @[main.scala 23:23]
  reg [7:0] fifo_83; // @[main.scala 23:23]
  reg [7:0] fifo_84; // @[main.scala 23:23]
  reg [7:0] fifo_85; // @[main.scala 23:23]
  reg [7:0] fifo_86; // @[main.scala 23:23]
  reg [7:0] fifo_87; // @[main.scala 23:23]
  reg [7:0] fifo_88; // @[main.scala 23:23]
  reg [7:0] fifo_89; // @[main.scala 23:23]
  reg [7:0] fifo_90; // @[main.scala 23:23]
  reg [7:0] fifo_91; // @[main.scala 23:23]
  reg [7:0] fifo_92; // @[main.scala 23:23]
  reg [7:0] fifo_93; // @[main.scala 23:23]
  reg [7:0] fifo_94; // @[main.scala 23:23]
  reg [7:0] fifo_95; // @[main.scala 23:23]
  reg [7:0] fifo_96; // @[main.scala 23:23]
  reg [7:0] fifo_97; // @[main.scala 23:23]
  reg [7:0] fifo_98; // @[main.scala 23:23]
  reg [7:0] fifo_99; // @[main.scala 23:23]
  reg [7:0] fifo_100; // @[main.scala 23:23]
  reg [7:0] fifo_101; // @[main.scala 23:23]
  reg [7:0] fifo_102; // @[main.scala 23:23]
  reg [7:0] fifo_103; // @[main.scala 23:23]
  reg [7:0] fifo_104; // @[main.scala 23:23]
  reg [7:0] fifo_105; // @[main.scala 23:23]
  reg [7:0] fifo_106; // @[main.scala 23:23]
  reg [7:0] fifo_107; // @[main.scala 23:23]
  reg [7:0] fifo_108; // @[main.scala 23:23]
  reg [7:0] fifo_109; // @[main.scala 23:23]
  reg [7:0] fifo_110; // @[main.scala 23:23]
  reg [7:0] fifo_111; // @[main.scala 23:23]
  reg [7:0] fifo_112; // @[main.scala 23:23]
  reg [7:0] fifo_113; // @[main.scala 23:23]
  reg [7:0] fifo_114; // @[main.scala 23:23]
  reg [7:0] fifo_115; // @[main.scala 23:23]
  reg [7:0] fifo_116; // @[main.scala 23:23]
  reg [7:0] fifo_117; // @[main.scala 23:23]
  reg [7:0] fifo_118; // @[main.scala 23:23]
  reg [7:0] fifo_119; // @[main.scala 23:23]
  reg [7:0] fifo_120; // @[main.scala 23:23]
  reg [7:0] fifo_121; // @[main.scala 23:23]
  reg [7:0] fifo_122; // @[main.scala 23:23]
  reg [7:0] fifo_123; // @[main.scala 23:23]
  reg [7:0] fifo_124; // @[main.scala 23:23]
  reg [7:0] fifo_125; // @[main.scala 23:23]
  reg [7:0] fifo_126; // @[main.scala 23:23]
  reg [7:0] fifo_127; // @[main.scala 23:23]
  reg [7:0] fifo_128; // @[main.scala 23:23]
  reg [7:0] fifo_129; // @[main.scala 23:23]
  reg [7:0] fifo_130; // @[main.scala 23:23]
  reg [7:0] fifo_131; // @[main.scala 23:23]
  reg [7:0] fifo_132; // @[main.scala 23:23]
  reg [7:0] fifo_133; // @[main.scala 23:23]
  reg [7:0] fifo_134; // @[main.scala 23:23]
  reg [7:0] fifo_135; // @[main.scala 23:23]
  reg [7:0] fifo_136; // @[main.scala 23:23]
  reg [7:0] fifo_137; // @[main.scala 23:23]
  reg [7:0] fifo_138; // @[main.scala 23:23]
  reg [7:0] fifo_139; // @[main.scala 23:23]
  reg [7:0] fifo_140; // @[main.scala 23:23]
  reg [7:0] fifo_141; // @[main.scala 23:23]
  reg [7:0] fifo_142; // @[main.scala 23:23]
  reg [7:0] fifo_143; // @[main.scala 23:23]
  reg [7:0] fifo_144; // @[main.scala 23:23]
  reg [7:0] fifo_145; // @[main.scala 23:23]
  reg [7:0] fifo_146; // @[main.scala 23:23]
  reg [7:0] fifo_147; // @[main.scala 23:23]
  reg [7:0] fifo_148; // @[main.scala 23:23]
  reg [7:0] fifo_149; // @[main.scala 23:23]
  reg [7:0] fifo_150; // @[main.scala 23:23]
  reg [7:0] fifo_151; // @[main.scala 23:23]
  reg [7:0] fifo_152; // @[main.scala 23:23]
  reg [7:0] fifo_153; // @[main.scala 23:23]
  reg [7:0] fifo_154; // @[main.scala 23:23]
  reg [7:0] fifo_155; // @[main.scala 23:23]
  reg [7:0] fifo_156; // @[main.scala 23:23]
  reg [7:0] fifo_157; // @[main.scala 23:23]
  reg [7:0] fifo_158; // @[main.scala 23:23]
  reg [7:0] fifo_159; // @[main.scala 23:23]
  reg [7:0] fifo_160; // @[main.scala 23:23]
  reg [7:0] fifo_161; // @[main.scala 23:23]
  reg [7:0] fifo_162; // @[main.scala 23:23]
  reg [7:0] fifo_163; // @[main.scala 23:23]
  reg [7:0] fifo_164; // @[main.scala 23:23]
  reg [7:0] fifo_165; // @[main.scala 23:23]
  reg [7:0] fifo_166; // @[main.scala 23:23]
  reg [7:0] fifo_167; // @[main.scala 23:23]
  reg [7:0] fifo_168; // @[main.scala 23:23]
  reg [7:0] fifo_169; // @[main.scala 23:23]
  reg [7:0] fifo_170; // @[main.scala 23:23]
  reg [7:0] fifo_171; // @[main.scala 23:23]
  reg [7:0] fifo_172; // @[main.scala 23:23]
  reg [7:0] fifo_173; // @[main.scala 23:23]
  reg [7:0] fifo_174; // @[main.scala 23:23]
  reg [7:0] fifo_175; // @[main.scala 23:23]
  reg [7:0] fifo_176; // @[main.scala 23:23]
  reg [7:0] fifo_177; // @[main.scala 23:23]
  reg [7:0] fifo_178; // @[main.scala 23:23]
  reg [7:0] fifo_179; // @[main.scala 23:23]
  reg [7:0] fifo_180; // @[main.scala 23:23]
  reg [7:0] fifo_181; // @[main.scala 23:23]
  reg [7:0] fifo_182; // @[main.scala 23:23]
  reg [7:0] fifo_183; // @[main.scala 23:23]
  reg [7:0] fifo_184; // @[main.scala 23:23]
  reg [7:0] fifo_185; // @[main.scala 23:23]
  reg [7:0] fifo_186; // @[main.scala 23:23]
  reg [7:0] fifo_187; // @[main.scala 23:23]
  reg [7:0] fifo_188; // @[main.scala 23:23]
  reg [7:0] fifo_189; // @[main.scala 23:23]
  reg [7:0] fifo_190; // @[main.scala 23:23]
  reg [7:0] fifo_191; // @[main.scala 23:23]
  reg [7:0] fifo_192; // @[main.scala 23:23]
  reg [7:0] fifo_193; // @[main.scala 23:23]
  reg [7:0] fifo_194; // @[main.scala 23:23]
  reg [7:0] fifo_195; // @[main.scala 23:23]
  reg [7:0] fifo_196; // @[main.scala 23:23]
  reg [7:0] fifo_197; // @[main.scala 23:23]
  reg [7:0] fifo_198; // @[main.scala 23:23]
  reg [7:0] fifo_199; // @[main.scala 23:23]
  reg [7:0] fifo_200; // @[main.scala 23:23]
  reg [7:0] fifo_201; // @[main.scala 23:23]
  reg [7:0] fifo_202; // @[main.scala 23:23]
  reg [7:0] fifo_203; // @[main.scala 23:23]
  reg [7:0] fifo_204; // @[main.scala 23:23]
  reg [7:0] fifo_205; // @[main.scala 23:23]
  reg [7:0] fifo_206; // @[main.scala 23:23]
  reg [7:0] fifo_207; // @[main.scala 23:23]
  reg [7:0] fifo_208; // @[main.scala 23:23]
  reg [7:0] fifo_209; // @[main.scala 23:23]
  reg [7:0] fifo_210; // @[main.scala 23:23]
  reg [7:0] fifo_211; // @[main.scala 23:23]
  reg [7:0] fifo_212; // @[main.scala 23:23]
  reg [7:0] fifo_213; // @[main.scala 23:23]
  reg [7:0] fifo_214; // @[main.scala 23:23]
  reg [7:0] fifo_215; // @[main.scala 23:23]
  reg [7:0] fifo_216; // @[main.scala 23:23]
  reg [7:0] fifo_217; // @[main.scala 23:23]
  reg [7:0] fifo_218; // @[main.scala 23:23]
  reg [7:0] fifo_219; // @[main.scala 23:23]
  reg [7:0] fifo_220; // @[main.scala 23:23]
  reg [7:0] fifo_221; // @[main.scala 23:23]
  reg [7:0] fifo_222; // @[main.scala 23:23]
  reg [7:0] fifo_223; // @[main.scala 23:23]
  reg [7:0] fifo_224; // @[main.scala 23:23]
  reg [7:0] fifo_225; // @[main.scala 23:23]
  reg [7:0] fifo_226; // @[main.scala 23:23]
  reg [7:0] fifo_227; // @[main.scala 23:23]
  reg [7:0] fifo_228; // @[main.scala 23:23]
  reg [7:0] fifo_229; // @[main.scala 23:23]
  reg [7:0] fifo_230; // @[main.scala 23:23]
  reg [7:0] fifo_231; // @[main.scala 23:23]
  reg [7:0] fifo_232; // @[main.scala 23:23]
  reg [7:0] fifo_233; // @[main.scala 23:23]
  reg [7:0] fifo_234; // @[main.scala 23:23]
  reg [7:0] fifo_235; // @[main.scala 23:23]
  reg [7:0] fifo_236; // @[main.scala 23:23]
  reg [7:0] fifo_237; // @[main.scala 23:23]
  reg [7:0] fifo_238; // @[main.scala 23:23]
  reg [7:0] fifo_239; // @[main.scala 23:23]
  reg [7:0] fifo_240; // @[main.scala 23:23]
  reg [7:0] fifo_241; // @[main.scala 23:23]
  reg [7:0] fifo_242; // @[main.scala 23:23]
  reg [7:0] fifo_243; // @[main.scala 23:23]
  reg [7:0] fifo_244; // @[main.scala 23:23]
  reg [7:0] fifo_245; // @[main.scala 23:23]
  reg [7:0] fifo_246; // @[main.scala 23:23]
  reg [7:0] fifo_247; // @[main.scala 23:23]
  reg [7:0] fifo_248; // @[main.scala 23:23]
  reg [7:0] fifo_249; // @[main.scala 23:23]
  reg [7:0] fifo_250; // @[main.scala 23:23]
  reg [7:0] fifo_251; // @[main.scala 23:23]
  reg [7:0] fifo_252; // @[main.scala 23:23]
  reg [7:0] fifo_253; // @[main.scala 23:23]
  reg [7:0] fifo_254; // @[main.scala 23:23]
  reg [7:0] fifo_255; // @[main.scala 23:23]
  wire [7:0] _GEN_257 = 8'h1 == io_in_addr ? fifo_1 : fifo_0; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_258 = 8'h2 == io_in_addr ? fifo_2 : _GEN_257; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_259 = 8'h3 == io_in_addr ? fifo_3 : _GEN_258; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_260 = 8'h4 == io_in_addr ? fifo_4 : _GEN_259; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_261 = 8'h5 == io_in_addr ? fifo_5 : _GEN_260; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_262 = 8'h6 == io_in_addr ? fifo_6 : _GEN_261; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_263 = 8'h7 == io_in_addr ? fifo_7 : _GEN_262; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_264 = 8'h8 == io_in_addr ? fifo_8 : _GEN_263; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_265 = 8'h9 == io_in_addr ? fifo_9 : _GEN_264; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_266 = 8'ha == io_in_addr ? fifo_10 : _GEN_265; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_267 = 8'hb == io_in_addr ? fifo_11 : _GEN_266; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_268 = 8'hc == io_in_addr ? fifo_12 : _GEN_267; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_269 = 8'hd == io_in_addr ? fifo_13 : _GEN_268; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_270 = 8'he == io_in_addr ? fifo_14 : _GEN_269; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_271 = 8'hf == io_in_addr ? fifo_15 : _GEN_270; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_272 = 8'h10 == io_in_addr ? fifo_16 : _GEN_271; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_273 = 8'h11 == io_in_addr ? fifo_17 : _GEN_272; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_274 = 8'h12 == io_in_addr ? fifo_18 : _GEN_273; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_275 = 8'h13 == io_in_addr ? fifo_19 : _GEN_274; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_276 = 8'h14 == io_in_addr ? fifo_20 : _GEN_275; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_277 = 8'h15 == io_in_addr ? fifo_21 : _GEN_276; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_278 = 8'h16 == io_in_addr ? fifo_22 : _GEN_277; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_279 = 8'h17 == io_in_addr ? fifo_23 : _GEN_278; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_280 = 8'h18 == io_in_addr ? fifo_24 : _GEN_279; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_281 = 8'h19 == io_in_addr ? fifo_25 : _GEN_280; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_282 = 8'h1a == io_in_addr ? fifo_26 : _GEN_281; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_283 = 8'h1b == io_in_addr ? fifo_27 : _GEN_282; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_284 = 8'h1c == io_in_addr ? fifo_28 : _GEN_283; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_285 = 8'h1d == io_in_addr ? fifo_29 : _GEN_284; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_286 = 8'h1e == io_in_addr ? fifo_30 : _GEN_285; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_287 = 8'h1f == io_in_addr ? fifo_31 : _GEN_286; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_288 = 8'h20 == io_in_addr ? fifo_32 : _GEN_287; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_289 = 8'h21 == io_in_addr ? fifo_33 : _GEN_288; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_290 = 8'h22 == io_in_addr ? fifo_34 : _GEN_289; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_291 = 8'h23 == io_in_addr ? fifo_35 : _GEN_290; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_292 = 8'h24 == io_in_addr ? fifo_36 : _GEN_291; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_293 = 8'h25 == io_in_addr ? fifo_37 : _GEN_292; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_294 = 8'h26 == io_in_addr ? fifo_38 : _GEN_293; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_295 = 8'h27 == io_in_addr ? fifo_39 : _GEN_294; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_296 = 8'h28 == io_in_addr ? fifo_40 : _GEN_295; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_297 = 8'h29 == io_in_addr ? fifo_41 : _GEN_296; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_298 = 8'h2a == io_in_addr ? fifo_42 : _GEN_297; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_299 = 8'h2b == io_in_addr ? fifo_43 : _GEN_298; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_300 = 8'h2c == io_in_addr ? fifo_44 : _GEN_299; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_301 = 8'h2d == io_in_addr ? fifo_45 : _GEN_300; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_302 = 8'h2e == io_in_addr ? fifo_46 : _GEN_301; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_303 = 8'h2f == io_in_addr ? fifo_47 : _GEN_302; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_304 = 8'h30 == io_in_addr ? fifo_48 : _GEN_303; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_305 = 8'h31 == io_in_addr ? fifo_49 : _GEN_304; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_306 = 8'h32 == io_in_addr ? fifo_50 : _GEN_305; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_307 = 8'h33 == io_in_addr ? fifo_51 : _GEN_306; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_308 = 8'h34 == io_in_addr ? fifo_52 : _GEN_307; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_309 = 8'h35 == io_in_addr ? fifo_53 : _GEN_308; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_310 = 8'h36 == io_in_addr ? fifo_54 : _GEN_309; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_311 = 8'h37 == io_in_addr ? fifo_55 : _GEN_310; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_312 = 8'h38 == io_in_addr ? fifo_56 : _GEN_311; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_313 = 8'h39 == io_in_addr ? fifo_57 : _GEN_312; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_314 = 8'h3a == io_in_addr ? fifo_58 : _GEN_313; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_315 = 8'h3b == io_in_addr ? fifo_59 : _GEN_314; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_316 = 8'h3c == io_in_addr ? fifo_60 : _GEN_315; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_317 = 8'h3d == io_in_addr ? fifo_61 : _GEN_316; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_318 = 8'h3e == io_in_addr ? fifo_62 : _GEN_317; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_319 = 8'h3f == io_in_addr ? fifo_63 : _GEN_318; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_320 = 8'h40 == io_in_addr ? fifo_64 : _GEN_319; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_321 = 8'h41 == io_in_addr ? fifo_65 : _GEN_320; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_322 = 8'h42 == io_in_addr ? fifo_66 : _GEN_321; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_323 = 8'h43 == io_in_addr ? fifo_67 : _GEN_322; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_324 = 8'h44 == io_in_addr ? fifo_68 : _GEN_323; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_325 = 8'h45 == io_in_addr ? fifo_69 : _GEN_324; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_326 = 8'h46 == io_in_addr ? fifo_70 : _GEN_325; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_327 = 8'h47 == io_in_addr ? fifo_71 : _GEN_326; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_328 = 8'h48 == io_in_addr ? fifo_72 : _GEN_327; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_329 = 8'h49 == io_in_addr ? fifo_73 : _GEN_328; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_330 = 8'h4a == io_in_addr ? fifo_74 : _GEN_329; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_331 = 8'h4b == io_in_addr ? fifo_75 : _GEN_330; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_332 = 8'h4c == io_in_addr ? fifo_76 : _GEN_331; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_333 = 8'h4d == io_in_addr ? fifo_77 : _GEN_332; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_334 = 8'h4e == io_in_addr ? fifo_78 : _GEN_333; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_335 = 8'h4f == io_in_addr ? fifo_79 : _GEN_334; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_336 = 8'h50 == io_in_addr ? fifo_80 : _GEN_335; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_337 = 8'h51 == io_in_addr ? fifo_81 : _GEN_336; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_338 = 8'h52 == io_in_addr ? fifo_82 : _GEN_337; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_339 = 8'h53 == io_in_addr ? fifo_83 : _GEN_338; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_340 = 8'h54 == io_in_addr ? fifo_84 : _GEN_339; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_341 = 8'h55 == io_in_addr ? fifo_85 : _GEN_340; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_342 = 8'h56 == io_in_addr ? fifo_86 : _GEN_341; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_343 = 8'h57 == io_in_addr ? fifo_87 : _GEN_342; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_344 = 8'h58 == io_in_addr ? fifo_88 : _GEN_343; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_345 = 8'h59 == io_in_addr ? fifo_89 : _GEN_344; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_346 = 8'h5a == io_in_addr ? fifo_90 : _GEN_345; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_347 = 8'h5b == io_in_addr ? fifo_91 : _GEN_346; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_348 = 8'h5c == io_in_addr ? fifo_92 : _GEN_347; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_349 = 8'h5d == io_in_addr ? fifo_93 : _GEN_348; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_350 = 8'h5e == io_in_addr ? fifo_94 : _GEN_349; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_351 = 8'h5f == io_in_addr ? fifo_95 : _GEN_350; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_352 = 8'h60 == io_in_addr ? fifo_96 : _GEN_351; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_353 = 8'h61 == io_in_addr ? fifo_97 : _GEN_352; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_354 = 8'h62 == io_in_addr ? fifo_98 : _GEN_353; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_355 = 8'h63 == io_in_addr ? fifo_99 : _GEN_354; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_356 = 8'h64 == io_in_addr ? fifo_100 : _GEN_355; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_357 = 8'h65 == io_in_addr ? fifo_101 : _GEN_356; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_358 = 8'h66 == io_in_addr ? fifo_102 : _GEN_357; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_359 = 8'h67 == io_in_addr ? fifo_103 : _GEN_358; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_360 = 8'h68 == io_in_addr ? fifo_104 : _GEN_359; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_361 = 8'h69 == io_in_addr ? fifo_105 : _GEN_360; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_362 = 8'h6a == io_in_addr ? fifo_106 : _GEN_361; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_363 = 8'h6b == io_in_addr ? fifo_107 : _GEN_362; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_364 = 8'h6c == io_in_addr ? fifo_108 : _GEN_363; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_365 = 8'h6d == io_in_addr ? fifo_109 : _GEN_364; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_366 = 8'h6e == io_in_addr ? fifo_110 : _GEN_365; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_367 = 8'h6f == io_in_addr ? fifo_111 : _GEN_366; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_368 = 8'h70 == io_in_addr ? fifo_112 : _GEN_367; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_369 = 8'h71 == io_in_addr ? fifo_113 : _GEN_368; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_370 = 8'h72 == io_in_addr ? fifo_114 : _GEN_369; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_371 = 8'h73 == io_in_addr ? fifo_115 : _GEN_370; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_372 = 8'h74 == io_in_addr ? fifo_116 : _GEN_371; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_373 = 8'h75 == io_in_addr ? fifo_117 : _GEN_372; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_374 = 8'h76 == io_in_addr ? fifo_118 : _GEN_373; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_375 = 8'h77 == io_in_addr ? fifo_119 : _GEN_374; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_376 = 8'h78 == io_in_addr ? fifo_120 : _GEN_375; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_377 = 8'h79 == io_in_addr ? fifo_121 : _GEN_376; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_378 = 8'h7a == io_in_addr ? fifo_122 : _GEN_377; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_379 = 8'h7b == io_in_addr ? fifo_123 : _GEN_378; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_380 = 8'h7c == io_in_addr ? fifo_124 : _GEN_379; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_381 = 8'h7d == io_in_addr ? fifo_125 : _GEN_380; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_382 = 8'h7e == io_in_addr ? fifo_126 : _GEN_381; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_383 = 8'h7f == io_in_addr ? fifo_127 : _GEN_382; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_384 = 8'h80 == io_in_addr ? fifo_128 : _GEN_383; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_385 = 8'h81 == io_in_addr ? fifo_129 : _GEN_384; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_386 = 8'h82 == io_in_addr ? fifo_130 : _GEN_385; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_387 = 8'h83 == io_in_addr ? fifo_131 : _GEN_386; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_388 = 8'h84 == io_in_addr ? fifo_132 : _GEN_387; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_389 = 8'h85 == io_in_addr ? fifo_133 : _GEN_388; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_390 = 8'h86 == io_in_addr ? fifo_134 : _GEN_389; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_391 = 8'h87 == io_in_addr ? fifo_135 : _GEN_390; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_392 = 8'h88 == io_in_addr ? fifo_136 : _GEN_391; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_393 = 8'h89 == io_in_addr ? fifo_137 : _GEN_392; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_394 = 8'h8a == io_in_addr ? fifo_138 : _GEN_393; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_395 = 8'h8b == io_in_addr ? fifo_139 : _GEN_394; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_396 = 8'h8c == io_in_addr ? fifo_140 : _GEN_395; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_397 = 8'h8d == io_in_addr ? fifo_141 : _GEN_396; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_398 = 8'h8e == io_in_addr ? fifo_142 : _GEN_397; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_399 = 8'h8f == io_in_addr ? fifo_143 : _GEN_398; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_400 = 8'h90 == io_in_addr ? fifo_144 : _GEN_399; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_401 = 8'h91 == io_in_addr ? fifo_145 : _GEN_400; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_402 = 8'h92 == io_in_addr ? fifo_146 : _GEN_401; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_403 = 8'h93 == io_in_addr ? fifo_147 : _GEN_402; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_404 = 8'h94 == io_in_addr ? fifo_148 : _GEN_403; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_405 = 8'h95 == io_in_addr ? fifo_149 : _GEN_404; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_406 = 8'h96 == io_in_addr ? fifo_150 : _GEN_405; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_407 = 8'h97 == io_in_addr ? fifo_151 : _GEN_406; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_408 = 8'h98 == io_in_addr ? fifo_152 : _GEN_407; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_409 = 8'h99 == io_in_addr ? fifo_153 : _GEN_408; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_410 = 8'h9a == io_in_addr ? fifo_154 : _GEN_409; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_411 = 8'h9b == io_in_addr ? fifo_155 : _GEN_410; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_412 = 8'h9c == io_in_addr ? fifo_156 : _GEN_411; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_413 = 8'h9d == io_in_addr ? fifo_157 : _GEN_412; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_414 = 8'h9e == io_in_addr ? fifo_158 : _GEN_413; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_415 = 8'h9f == io_in_addr ? fifo_159 : _GEN_414; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_416 = 8'ha0 == io_in_addr ? fifo_160 : _GEN_415; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_417 = 8'ha1 == io_in_addr ? fifo_161 : _GEN_416; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_418 = 8'ha2 == io_in_addr ? fifo_162 : _GEN_417; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_419 = 8'ha3 == io_in_addr ? fifo_163 : _GEN_418; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_420 = 8'ha4 == io_in_addr ? fifo_164 : _GEN_419; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_421 = 8'ha5 == io_in_addr ? fifo_165 : _GEN_420; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_422 = 8'ha6 == io_in_addr ? fifo_166 : _GEN_421; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_423 = 8'ha7 == io_in_addr ? fifo_167 : _GEN_422; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_424 = 8'ha8 == io_in_addr ? fifo_168 : _GEN_423; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_425 = 8'ha9 == io_in_addr ? fifo_169 : _GEN_424; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_426 = 8'haa == io_in_addr ? fifo_170 : _GEN_425; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_427 = 8'hab == io_in_addr ? fifo_171 : _GEN_426; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_428 = 8'hac == io_in_addr ? fifo_172 : _GEN_427; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_429 = 8'had == io_in_addr ? fifo_173 : _GEN_428; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_430 = 8'hae == io_in_addr ? fifo_174 : _GEN_429; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_431 = 8'haf == io_in_addr ? fifo_175 : _GEN_430; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_432 = 8'hb0 == io_in_addr ? fifo_176 : _GEN_431; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_433 = 8'hb1 == io_in_addr ? fifo_177 : _GEN_432; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_434 = 8'hb2 == io_in_addr ? fifo_178 : _GEN_433; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_435 = 8'hb3 == io_in_addr ? fifo_179 : _GEN_434; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_436 = 8'hb4 == io_in_addr ? fifo_180 : _GEN_435; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_437 = 8'hb5 == io_in_addr ? fifo_181 : _GEN_436; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_438 = 8'hb6 == io_in_addr ? fifo_182 : _GEN_437; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_439 = 8'hb7 == io_in_addr ? fifo_183 : _GEN_438; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_440 = 8'hb8 == io_in_addr ? fifo_184 : _GEN_439; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_441 = 8'hb9 == io_in_addr ? fifo_185 : _GEN_440; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_442 = 8'hba == io_in_addr ? fifo_186 : _GEN_441; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_443 = 8'hbb == io_in_addr ? fifo_187 : _GEN_442; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_444 = 8'hbc == io_in_addr ? fifo_188 : _GEN_443; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_445 = 8'hbd == io_in_addr ? fifo_189 : _GEN_444; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_446 = 8'hbe == io_in_addr ? fifo_190 : _GEN_445; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_447 = 8'hbf == io_in_addr ? fifo_191 : _GEN_446; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_448 = 8'hc0 == io_in_addr ? fifo_192 : _GEN_447; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_449 = 8'hc1 == io_in_addr ? fifo_193 : _GEN_448; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_450 = 8'hc2 == io_in_addr ? fifo_194 : _GEN_449; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_451 = 8'hc3 == io_in_addr ? fifo_195 : _GEN_450; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_452 = 8'hc4 == io_in_addr ? fifo_196 : _GEN_451; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_453 = 8'hc5 == io_in_addr ? fifo_197 : _GEN_452; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_454 = 8'hc6 == io_in_addr ? fifo_198 : _GEN_453; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_455 = 8'hc7 == io_in_addr ? fifo_199 : _GEN_454; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_456 = 8'hc8 == io_in_addr ? fifo_200 : _GEN_455; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_457 = 8'hc9 == io_in_addr ? fifo_201 : _GEN_456; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_458 = 8'hca == io_in_addr ? fifo_202 : _GEN_457; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_459 = 8'hcb == io_in_addr ? fifo_203 : _GEN_458; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_460 = 8'hcc == io_in_addr ? fifo_204 : _GEN_459; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_461 = 8'hcd == io_in_addr ? fifo_205 : _GEN_460; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_462 = 8'hce == io_in_addr ? fifo_206 : _GEN_461; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_463 = 8'hcf == io_in_addr ? fifo_207 : _GEN_462; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_464 = 8'hd0 == io_in_addr ? fifo_208 : _GEN_463; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_465 = 8'hd1 == io_in_addr ? fifo_209 : _GEN_464; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_466 = 8'hd2 == io_in_addr ? fifo_210 : _GEN_465; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_467 = 8'hd3 == io_in_addr ? fifo_211 : _GEN_466; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_468 = 8'hd4 == io_in_addr ? fifo_212 : _GEN_467; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_469 = 8'hd5 == io_in_addr ? fifo_213 : _GEN_468; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_470 = 8'hd6 == io_in_addr ? fifo_214 : _GEN_469; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_471 = 8'hd7 == io_in_addr ? fifo_215 : _GEN_470; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_472 = 8'hd8 == io_in_addr ? fifo_216 : _GEN_471; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_473 = 8'hd9 == io_in_addr ? fifo_217 : _GEN_472; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_474 = 8'hda == io_in_addr ? fifo_218 : _GEN_473; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_475 = 8'hdb == io_in_addr ? fifo_219 : _GEN_474; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_476 = 8'hdc == io_in_addr ? fifo_220 : _GEN_475; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_477 = 8'hdd == io_in_addr ? fifo_221 : _GEN_476; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_478 = 8'hde == io_in_addr ? fifo_222 : _GEN_477; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_479 = 8'hdf == io_in_addr ? fifo_223 : _GEN_478; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_480 = 8'he0 == io_in_addr ? fifo_224 : _GEN_479; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_481 = 8'he1 == io_in_addr ? fifo_225 : _GEN_480; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_482 = 8'he2 == io_in_addr ? fifo_226 : _GEN_481; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_483 = 8'he3 == io_in_addr ? fifo_227 : _GEN_482; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_484 = 8'he4 == io_in_addr ? fifo_228 : _GEN_483; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_485 = 8'he5 == io_in_addr ? fifo_229 : _GEN_484; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_486 = 8'he6 == io_in_addr ? fifo_230 : _GEN_485; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_487 = 8'he7 == io_in_addr ? fifo_231 : _GEN_486; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_488 = 8'he8 == io_in_addr ? fifo_232 : _GEN_487; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_489 = 8'he9 == io_in_addr ? fifo_233 : _GEN_488; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_490 = 8'hea == io_in_addr ? fifo_234 : _GEN_489; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_491 = 8'heb == io_in_addr ? fifo_235 : _GEN_490; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_492 = 8'hec == io_in_addr ? fifo_236 : _GEN_491; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_493 = 8'hed == io_in_addr ? fifo_237 : _GEN_492; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_494 = 8'hee == io_in_addr ? fifo_238 : _GEN_493; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_495 = 8'hef == io_in_addr ? fifo_239 : _GEN_494; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_496 = 8'hf0 == io_in_addr ? fifo_240 : _GEN_495; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_497 = 8'hf1 == io_in_addr ? fifo_241 : _GEN_496; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_498 = 8'hf2 == io_in_addr ? fifo_242 : _GEN_497; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_499 = 8'hf3 == io_in_addr ? fifo_243 : _GEN_498; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_500 = 8'hf4 == io_in_addr ? fifo_244 : _GEN_499; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_501 = 8'hf5 == io_in_addr ? fifo_245 : _GEN_500; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_502 = 8'hf6 == io_in_addr ? fifo_246 : _GEN_501; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_503 = 8'hf7 == io_in_addr ? fifo_247 : _GEN_502; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_504 = 8'hf8 == io_in_addr ? fifo_248 : _GEN_503; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_505 = 8'hf9 == io_in_addr ? fifo_249 : _GEN_504; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_506 = 8'hfa == io_in_addr ? fifo_250 : _GEN_505; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_507 = 8'hfb == io_in_addr ? fifo_251 : _GEN_506; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_508 = 8'hfc == io_in_addr ? fifo_252 : _GEN_507; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_509 = 8'hfd == io_in_addr ? fifo_253 : _GEN_508; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_510 = 8'hfe == io_in_addr ? fifo_254 : _GEN_509; // @[main.scala 34:{21,21}]
  wire [7:0] _GEN_511 = 8'hff == io_in_addr ? fifo_255 : _GEN_510; // @[main.scala 34:{21,21}]
  assign io_out_data = io_in_en ? 8'h0 : _GEN_511; // @[main.scala 26:21 30:21 34:21]
  assign io_out_en = io_in_en ? 1'h0 : 1'h1; // @[main.scala 26:21 29:19 35:19]
  always @(posedge clock) begin
    if (reset) begin // @[main.scala 23:23]
      fifo_0 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h0 == io_in_addr) begin // @[main.scala 28:26]
        fifo_0 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_1 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h1 == io_in_addr) begin // @[main.scala 28:26]
        fifo_1 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_2 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h2 == io_in_addr) begin // @[main.scala 28:26]
        fifo_2 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_3 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h3 == io_in_addr) begin // @[main.scala 28:26]
        fifo_3 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_4 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h4 == io_in_addr) begin // @[main.scala 28:26]
        fifo_4 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_5 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h5 == io_in_addr) begin // @[main.scala 28:26]
        fifo_5 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_6 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h6 == io_in_addr) begin // @[main.scala 28:26]
        fifo_6 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_7 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h7 == io_in_addr) begin // @[main.scala 28:26]
        fifo_7 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_8 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h8 == io_in_addr) begin // @[main.scala 28:26]
        fifo_8 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_9 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h9 == io_in_addr) begin // @[main.scala 28:26]
        fifo_9 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_10 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha == io_in_addr) begin // @[main.scala 28:26]
        fifo_10 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_11 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb == io_in_addr) begin // @[main.scala 28:26]
        fifo_11 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_12 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc == io_in_addr) begin // @[main.scala 28:26]
        fifo_12 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_13 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd == io_in_addr) begin // @[main.scala 28:26]
        fifo_13 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_14 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he == io_in_addr) begin // @[main.scala 28:26]
        fifo_14 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_15 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf == io_in_addr) begin // @[main.scala 28:26]
        fifo_15 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_16 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h10 == io_in_addr) begin // @[main.scala 28:26]
        fifo_16 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_17 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h11 == io_in_addr) begin // @[main.scala 28:26]
        fifo_17 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_18 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h12 == io_in_addr) begin // @[main.scala 28:26]
        fifo_18 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_19 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h13 == io_in_addr) begin // @[main.scala 28:26]
        fifo_19 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_20 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h14 == io_in_addr) begin // @[main.scala 28:26]
        fifo_20 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_21 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h15 == io_in_addr) begin // @[main.scala 28:26]
        fifo_21 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_22 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h16 == io_in_addr) begin // @[main.scala 28:26]
        fifo_22 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_23 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h17 == io_in_addr) begin // @[main.scala 28:26]
        fifo_23 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_24 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h18 == io_in_addr) begin // @[main.scala 28:26]
        fifo_24 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_25 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h19 == io_in_addr) begin // @[main.scala 28:26]
        fifo_25 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_26 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h1a == io_in_addr) begin // @[main.scala 28:26]
        fifo_26 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_27 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h1b == io_in_addr) begin // @[main.scala 28:26]
        fifo_27 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_28 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h1c == io_in_addr) begin // @[main.scala 28:26]
        fifo_28 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_29 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h1d == io_in_addr) begin // @[main.scala 28:26]
        fifo_29 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_30 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h1e == io_in_addr) begin // @[main.scala 28:26]
        fifo_30 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_31 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h1f == io_in_addr) begin // @[main.scala 28:26]
        fifo_31 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_32 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h20 == io_in_addr) begin // @[main.scala 28:26]
        fifo_32 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_33 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h21 == io_in_addr) begin // @[main.scala 28:26]
        fifo_33 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_34 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h22 == io_in_addr) begin // @[main.scala 28:26]
        fifo_34 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_35 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h23 == io_in_addr) begin // @[main.scala 28:26]
        fifo_35 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_36 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h24 == io_in_addr) begin // @[main.scala 28:26]
        fifo_36 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_37 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h25 == io_in_addr) begin // @[main.scala 28:26]
        fifo_37 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_38 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h26 == io_in_addr) begin // @[main.scala 28:26]
        fifo_38 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_39 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h27 == io_in_addr) begin // @[main.scala 28:26]
        fifo_39 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_40 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h28 == io_in_addr) begin // @[main.scala 28:26]
        fifo_40 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_41 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h29 == io_in_addr) begin // @[main.scala 28:26]
        fifo_41 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_42 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h2a == io_in_addr) begin // @[main.scala 28:26]
        fifo_42 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_43 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h2b == io_in_addr) begin // @[main.scala 28:26]
        fifo_43 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_44 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h2c == io_in_addr) begin // @[main.scala 28:26]
        fifo_44 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_45 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h2d == io_in_addr) begin // @[main.scala 28:26]
        fifo_45 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_46 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h2e == io_in_addr) begin // @[main.scala 28:26]
        fifo_46 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_47 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h2f == io_in_addr) begin // @[main.scala 28:26]
        fifo_47 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_48 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h30 == io_in_addr) begin // @[main.scala 28:26]
        fifo_48 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_49 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h31 == io_in_addr) begin // @[main.scala 28:26]
        fifo_49 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_50 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h32 == io_in_addr) begin // @[main.scala 28:26]
        fifo_50 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_51 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h33 == io_in_addr) begin // @[main.scala 28:26]
        fifo_51 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_52 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h34 == io_in_addr) begin // @[main.scala 28:26]
        fifo_52 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_53 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h35 == io_in_addr) begin // @[main.scala 28:26]
        fifo_53 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_54 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h36 == io_in_addr) begin // @[main.scala 28:26]
        fifo_54 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_55 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h37 == io_in_addr) begin // @[main.scala 28:26]
        fifo_55 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_56 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h38 == io_in_addr) begin // @[main.scala 28:26]
        fifo_56 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_57 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h39 == io_in_addr) begin // @[main.scala 28:26]
        fifo_57 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_58 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h3a == io_in_addr) begin // @[main.scala 28:26]
        fifo_58 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_59 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h3b == io_in_addr) begin // @[main.scala 28:26]
        fifo_59 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_60 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h3c == io_in_addr) begin // @[main.scala 28:26]
        fifo_60 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_61 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h3d == io_in_addr) begin // @[main.scala 28:26]
        fifo_61 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_62 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h3e == io_in_addr) begin // @[main.scala 28:26]
        fifo_62 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_63 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h3f == io_in_addr) begin // @[main.scala 28:26]
        fifo_63 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_64 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h40 == io_in_addr) begin // @[main.scala 28:26]
        fifo_64 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_65 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h41 == io_in_addr) begin // @[main.scala 28:26]
        fifo_65 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_66 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h42 == io_in_addr) begin // @[main.scala 28:26]
        fifo_66 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_67 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h43 == io_in_addr) begin // @[main.scala 28:26]
        fifo_67 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_68 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h44 == io_in_addr) begin // @[main.scala 28:26]
        fifo_68 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_69 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h45 == io_in_addr) begin // @[main.scala 28:26]
        fifo_69 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_70 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h46 == io_in_addr) begin // @[main.scala 28:26]
        fifo_70 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_71 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h47 == io_in_addr) begin // @[main.scala 28:26]
        fifo_71 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_72 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h48 == io_in_addr) begin // @[main.scala 28:26]
        fifo_72 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_73 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h49 == io_in_addr) begin // @[main.scala 28:26]
        fifo_73 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_74 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h4a == io_in_addr) begin // @[main.scala 28:26]
        fifo_74 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_75 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h4b == io_in_addr) begin // @[main.scala 28:26]
        fifo_75 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_76 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h4c == io_in_addr) begin // @[main.scala 28:26]
        fifo_76 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_77 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h4d == io_in_addr) begin // @[main.scala 28:26]
        fifo_77 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_78 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h4e == io_in_addr) begin // @[main.scala 28:26]
        fifo_78 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_79 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h4f == io_in_addr) begin // @[main.scala 28:26]
        fifo_79 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_80 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h50 == io_in_addr) begin // @[main.scala 28:26]
        fifo_80 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_81 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h51 == io_in_addr) begin // @[main.scala 28:26]
        fifo_81 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_82 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h52 == io_in_addr) begin // @[main.scala 28:26]
        fifo_82 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_83 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h53 == io_in_addr) begin // @[main.scala 28:26]
        fifo_83 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_84 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h54 == io_in_addr) begin // @[main.scala 28:26]
        fifo_84 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_85 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h55 == io_in_addr) begin // @[main.scala 28:26]
        fifo_85 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_86 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h56 == io_in_addr) begin // @[main.scala 28:26]
        fifo_86 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_87 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h57 == io_in_addr) begin // @[main.scala 28:26]
        fifo_87 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_88 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h58 == io_in_addr) begin // @[main.scala 28:26]
        fifo_88 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_89 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h59 == io_in_addr) begin // @[main.scala 28:26]
        fifo_89 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_90 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h5a == io_in_addr) begin // @[main.scala 28:26]
        fifo_90 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_91 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h5b == io_in_addr) begin // @[main.scala 28:26]
        fifo_91 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_92 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h5c == io_in_addr) begin // @[main.scala 28:26]
        fifo_92 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_93 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h5d == io_in_addr) begin // @[main.scala 28:26]
        fifo_93 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_94 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h5e == io_in_addr) begin // @[main.scala 28:26]
        fifo_94 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_95 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h5f == io_in_addr) begin // @[main.scala 28:26]
        fifo_95 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_96 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h60 == io_in_addr) begin // @[main.scala 28:26]
        fifo_96 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_97 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h61 == io_in_addr) begin // @[main.scala 28:26]
        fifo_97 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_98 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h62 == io_in_addr) begin // @[main.scala 28:26]
        fifo_98 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_99 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h63 == io_in_addr) begin // @[main.scala 28:26]
        fifo_99 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_100 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h64 == io_in_addr) begin // @[main.scala 28:26]
        fifo_100 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_101 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h65 == io_in_addr) begin // @[main.scala 28:26]
        fifo_101 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_102 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h66 == io_in_addr) begin // @[main.scala 28:26]
        fifo_102 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_103 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h67 == io_in_addr) begin // @[main.scala 28:26]
        fifo_103 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_104 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h68 == io_in_addr) begin // @[main.scala 28:26]
        fifo_104 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_105 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h69 == io_in_addr) begin // @[main.scala 28:26]
        fifo_105 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_106 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h6a == io_in_addr) begin // @[main.scala 28:26]
        fifo_106 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_107 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h6b == io_in_addr) begin // @[main.scala 28:26]
        fifo_107 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_108 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h6c == io_in_addr) begin // @[main.scala 28:26]
        fifo_108 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_109 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h6d == io_in_addr) begin // @[main.scala 28:26]
        fifo_109 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_110 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h6e == io_in_addr) begin // @[main.scala 28:26]
        fifo_110 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_111 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h6f == io_in_addr) begin // @[main.scala 28:26]
        fifo_111 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_112 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h70 == io_in_addr) begin // @[main.scala 28:26]
        fifo_112 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_113 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h71 == io_in_addr) begin // @[main.scala 28:26]
        fifo_113 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_114 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h72 == io_in_addr) begin // @[main.scala 28:26]
        fifo_114 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_115 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h73 == io_in_addr) begin // @[main.scala 28:26]
        fifo_115 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_116 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h74 == io_in_addr) begin // @[main.scala 28:26]
        fifo_116 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_117 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h75 == io_in_addr) begin // @[main.scala 28:26]
        fifo_117 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_118 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h76 == io_in_addr) begin // @[main.scala 28:26]
        fifo_118 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_119 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h77 == io_in_addr) begin // @[main.scala 28:26]
        fifo_119 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_120 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h78 == io_in_addr) begin // @[main.scala 28:26]
        fifo_120 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_121 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h79 == io_in_addr) begin // @[main.scala 28:26]
        fifo_121 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_122 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h7a == io_in_addr) begin // @[main.scala 28:26]
        fifo_122 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_123 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h7b == io_in_addr) begin // @[main.scala 28:26]
        fifo_123 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_124 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h7c == io_in_addr) begin // @[main.scala 28:26]
        fifo_124 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_125 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h7d == io_in_addr) begin // @[main.scala 28:26]
        fifo_125 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_126 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h7e == io_in_addr) begin // @[main.scala 28:26]
        fifo_126 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_127 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h7f == io_in_addr) begin // @[main.scala 28:26]
        fifo_127 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_128 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h80 == io_in_addr) begin // @[main.scala 28:26]
        fifo_128 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_129 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h81 == io_in_addr) begin // @[main.scala 28:26]
        fifo_129 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_130 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h82 == io_in_addr) begin // @[main.scala 28:26]
        fifo_130 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_131 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h83 == io_in_addr) begin // @[main.scala 28:26]
        fifo_131 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_132 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h84 == io_in_addr) begin // @[main.scala 28:26]
        fifo_132 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_133 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h85 == io_in_addr) begin // @[main.scala 28:26]
        fifo_133 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_134 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h86 == io_in_addr) begin // @[main.scala 28:26]
        fifo_134 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_135 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h87 == io_in_addr) begin // @[main.scala 28:26]
        fifo_135 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_136 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h88 == io_in_addr) begin // @[main.scala 28:26]
        fifo_136 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_137 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h89 == io_in_addr) begin // @[main.scala 28:26]
        fifo_137 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_138 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h8a == io_in_addr) begin // @[main.scala 28:26]
        fifo_138 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_139 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h8b == io_in_addr) begin // @[main.scala 28:26]
        fifo_139 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_140 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h8c == io_in_addr) begin // @[main.scala 28:26]
        fifo_140 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_141 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h8d == io_in_addr) begin // @[main.scala 28:26]
        fifo_141 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_142 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h8e == io_in_addr) begin // @[main.scala 28:26]
        fifo_142 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_143 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h8f == io_in_addr) begin // @[main.scala 28:26]
        fifo_143 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_144 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h90 == io_in_addr) begin // @[main.scala 28:26]
        fifo_144 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_145 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h91 == io_in_addr) begin // @[main.scala 28:26]
        fifo_145 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_146 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h92 == io_in_addr) begin // @[main.scala 28:26]
        fifo_146 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_147 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h93 == io_in_addr) begin // @[main.scala 28:26]
        fifo_147 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_148 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h94 == io_in_addr) begin // @[main.scala 28:26]
        fifo_148 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_149 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h95 == io_in_addr) begin // @[main.scala 28:26]
        fifo_149 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_150 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h96 == io_in_addr) begin // @[main.scala 28:26]
        fifo_150 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_151 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h97 == io_in_addr) begin // @[main.scala 28:26]
        fifo_151 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_152 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h98 == io_in_addr) begin // @[main.scala 28:26]
        fifo_152 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_153 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h99 == io_in_addr) begin // @[main.scala 28:26]
        fifo_153 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_154 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h9a == io_in_addr) begin // @[main.scala 28:26]
        fifo_154 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_155 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h9b == io_in_addr) begin // @[main.scala 28:26]
        fifo_155 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_156 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h9c == io_in_addr) begin // @[main.scala 28:26]
        fifo_156 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_157 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h9d == io_in_addr) begin // @[main.scala 28:26]
        fifo_157 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_158 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h9e == io_in_addr) begin // @[main.scala 28:26]
        fifo_158 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_159 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'h9f == io_in_addr) begin // @[main.scala 28:26]
        fifo_159 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_160 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha0 == io_in_addr) begin // @[main.scala 28:26]
        fifo_160 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_161 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha1 == io_in_addr) begin // @[main.scala 28:26]
        fifo_161 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_162 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha2 == io_in_addr) begin // @[main.scala 28:26]
        fifo_162 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_163 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha3 == io_in_addr) begin // @[main.scala 28:26]
        fifo_163 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_164 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha4 == io_in_addr) begin // @[main.scala 28:26]
        fifo_164 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_165 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha5 == io_in_addr) begin // @[main.scala 28:26]
        fifo_165 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_166 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha6 == io_in_addr) begin // @[main.scala 28:26]
        fifo_166 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_167 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha7 == io_in_addr) begin // @[main.scala 28:26]
        fifo_167 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_168 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha8 == io_in_addr) begin // @[main.scala 28:26]
        fifo_168 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_169 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'ha9 == io_in_addr) begin // @[main.scala 28:26]
        fifo_169 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_170 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'haa == io_in_addr) begin // @[main.scala 28:26]
        fifo_170 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_171 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hab == io_in_addr) begin // @[main.scala 28:26]
        fifo_171 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_172 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hac == io_in_addr) begin // @[main.scala 28:26]
        fifo_172 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_173 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'had == io_in_addr) begin // @[main.scala 28:26]
        fifo_173 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_174 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hae == io_in_addr) begin // @[main.scala 28:26]
        fifo_174 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_175 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'haf == io_in_addr) begin // @[main.scala 28:26]
        fifo_175 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_176 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb0 == io_in_addr) begin // @[main.scala 28:26]
        fifo_176 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_177 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb1 == io_in_addr) begin // @[main.scala 28:26]
        fifo_177 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_178 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb2 == io_in_addr) begin // @[main.scala 28:26]
        fifo_178 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_179 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb3 == io_in_addr) begin // @[main.scala 28:26]
        fifo_179 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_180 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb4 == io_in_addr) begin // @[main.scala 28:26]
        fifo_180 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_181 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb5 == io_in_addr) begin // @[main.scala 28:26]
        fifo_181 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_182 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb6 == io_in_addr) begin // @[main.scala 28:26]
        fifo_182 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_183 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb7 == io_in_addr) begin // @[main.scala 28:26]
        fifo_183 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_184 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb8 == io_in_addr) begin // @[main.scala 28:26]
        fifo_184 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_185 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hb9 == io_in_addr) begin // @[main.scala 28:26]
        fifo_185 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_186 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hba == io_in_addr) begin // @[main.scala 28:26]
        fifo_186 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_187 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hbb == io_in_addr) begin // @[main.scala 28:26]
        fifo_187 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_188 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hbc == io_in_addr) begin // @[main.scala 28:26]
        fifo_188 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_189 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hbd == io_in_addr) begin // @[main.scala 28:26]
        fifo_189 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_190 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hbe == io_in_addr) begin // @[main.scala 28:26]
        fifo_190 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_191 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hbf == io_in_addr) begin // @[main.scala 28:26]
        fifo_191 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_192 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc0 == io_in_addr) begin // @[main.scala 28:26]
        fifo_192 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_193 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc1 == io_in_addr) begin // @[main.scala 28:26]
        fifo_193 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_194 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc2 == io_in_addr) begin // @[main.scala 28:26]
        fifo_194 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_195 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc3 == io_in_addr) begin // @[main.scala 28:26]
        fifo_195 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_196 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc4 == io_in_addr) begin // @[main.scala 28:26]
        fifo_196 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_197 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc5 == io_in_addr) begin // @[main.scala 28:26]
        fifo_197 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_198 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc6 == io_in_addr) begin // @[main.scala 28:26]
        fifo_198 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_199 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc7 == io_in_addr) begin // @[main.scala 28:26]
        fifo_199 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_200 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc8 == io_in_addr) begin // @[main.scala 28:26]
        fifo_200 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_201 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hc9 == io_in_addr) begin // @[main.scala 28:26]
        fifo_201 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_202 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hca == io_in_addr) begin // @[main.scala 28:26]
        fifo_202 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_203 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hcb == io_in_addr) begin // @[main.scala 28:26]
        fifo_203 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_204 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hcc == io_in_addr) begin // @[main.scala 28:26]
        fifo_204 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_205 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hcd == io_in_addr) begin // @[main.scala 28:26]
        fifo_205 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_206 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hce == io_in_addr) begin // @[main.scala 28:26]
        fifo_206 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_207 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hcf == io_in_addr) begin // @[main.scala 28:26]
        fifo_207 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_208 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd0 == io_in_addr) begin // @[main.scala 28:26]
        fifo_208 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_209 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd1 == io_in_addr) begin // @[main.scala 28:26]
        fifo_209 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_210 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd2 == io_in_addr) begin // @[main.scala 28:26]
        fifo_210 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_211 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd3 == io_in_addr) begin // @[main.scala 28:26]
        fifo_211 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_212 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd4 == io_in_addr) begin // @[main.scala 28:26]
        fifo_212 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_213 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd5 == io_in_addr) begin // @[main.scala 28:26]
        fifo_213 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_214 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd6 == io_in_addr) begin // @[main.scala 28:26]
        fifo_214 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_215 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd7 == io_in_addr) begin // @[main.scala 28:26]
        fifo_215 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_216 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd8 == io_in_addr) begin // @[main.scala 28:26]
        fifo_216 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_217 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hd9 == io_in_addr) begin // @[main.scala 28:26]
        fifo_217 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_218 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hda == io_in_addr) begin // @[main.scala 28:26]
        fifo_218 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_219 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hdb == io_in_addr) begin // @[main.scala 28:26]
        fifo_219 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_220 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hdc == io_in_addr) begin // @[main.scala 28:26]
        fifo_220 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_221 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hdd == io_in_addr) begin // @[main.scala 28:26]
        fifo_221 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_222 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hde == io_in_addr) begin // @[main.scala 28:26]
        fifo_222 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_223 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hdf == io_in_addr) begin // @[main.scala 28:26]
        fifo_223 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_224 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he0 == io_in_addr) begin // @[main.scala 28:26]
        fifo_224 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_225 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he1 == io_in_addr) begin // @[main.scala 28:26]
        fifo_225 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_226 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he2 == io_in_addr) begin // @[main.scala 28:26]
        fifo_226 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_227 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he3 == io_in_addr) begin // @[main.scala 28:26]
        fifo_227 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_228 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he4 == io_in_addr) begin // @[main.scala 28:26]
        fifo_228 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_229 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he5 == io_in_addr) begin // @[main.scala 28:26]
        fifo_229 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_230 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he6 == io_in_addr) begin // @[main.scala 28:26]
        fifo_230 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_231 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he7 == io_in_addr) begin // @[main.scala 28:26]
        fifo_231 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_232 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he8 == io_in_addr) begin // @[main.scala 28:26]
        fifo_232 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_233 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'he9 == io_in_addr) begin // @[main.scala 28:26]
        fifo_233 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_234 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hea == io_in_addr) begin // @[main.scala 28:26]
        fifo_234 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_235 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'heb == io_in_addr) begin // @[main.scala 28:26]
        fifo_235 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_236 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hec == io_in_addr) begin // @[main.scala 28:26]
        fifo_236 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_237 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hed == io_in_addr) begin // @[main.scala 28:26]
        fifo_237 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_238 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hee == io_in_addr) begin // @[main.scala 28:26]
        fifo_238 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_239 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hef == io_in_addr) begin // @[main.scala 28:26]
        fifo_239 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_240 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf0 == io_in_addr) begin // @[main.scala 28:26]
        fifo_240 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_241 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf1 == io_in_addr) begin // @[main.scala 28:26]
        fifo_241 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_242 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf2 == io_in_addr) begin // @[main.scala 28:26]
        fifo_242 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_243 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf3 == io_in_addr) begin // @[main.scala 28:26]
        fifo_243 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_244 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf4 == io_in_addr) begin // @[main.scala 28:26]
        fifo_244 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_245 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf5 == io_in_addr) begin // @[main.scala 28:26]
        fifo_245 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_246 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf6 == io_in_addr) begin // @[main.scala 28:26]
        fifo_246 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_247 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf7 == io_in_addr) begin // @[main.scala 28:26]
        fifo_247 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_248 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf8 == io_in_addr) begin // @[main.scala 28:26]
        fifo_248 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_249 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hf9 == io_in_addr) begin // @[main.scala 28:26]
        fifo_249 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_250 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hfa == io_in_addr) begin // @[main.scala 28:26]
        fifo_250 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_251 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hfb == io_in_addr) begin // @[main.scala 28:26]
        fifo_251 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_252 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hfc == io_in_addr) begin // @[main.scala 28:26]
        fifo_252 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_253 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hfd == io_in_addr) begin // @[main.scala 28:26]
        fifo_253 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_254 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hfe == io_in_addr) begin // @[main.scala 28:26]
        fifo_254 <= io_in_data; // @[main.scala 28:26]
      end
    end
    if (reset) begin // @[main.scala 23:23]
      fifo_255 <= 8'h0; // @[main.scala 23:23]
    end else if (io_in_en) begin // @[main.scala 26:21]
      if (8'hff == io_in_addr) begin // @[main.scala 28:26]
        fifo_255 <= io_in_data; // @[main.scala 28:26]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fifo_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  fifo_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  fifo_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  fifo_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  fifo_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  fifo_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  fifo_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  fifo_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  fifo_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  fifo_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  fifo_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  fifo_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  fifo_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  fifo_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  fifo_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  fifo_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  fifo_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  fifo_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  fifo_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  fifo_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  fifo_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  fifo_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  fifo_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  fifo_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  fifo_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  fifo_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  fifo_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  fifo_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  fifo_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  fifo_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  fifo_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  fifo_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  fifo_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  fifo_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  fifo_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  fifo_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  fifo_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  fifo_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  fifo_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  fifo_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  fifo_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  fifo_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  fifo_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  fifo_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  fifo_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  fifo_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  fifo_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  fifo_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  fifo_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  fifo_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  fifo_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  fifo_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  fifo_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  fifo_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  fifo_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  fifo_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  fifo_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  fifo_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  fifo_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  fifo_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  fifo_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  fifo_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  fifo_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  fifo_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  fifo_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  fifo_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  fifo_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  fifo_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  fifo_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  fifo_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  fifo_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  fifo_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  fifo_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  fifo_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  fifo_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  fifo_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  fifo_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  fifo_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  fifo_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  fifo_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  fifo_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  fifo_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  fifo_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  fifo_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  fifo_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  fifo_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  fifo_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  fifo_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  fifo_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  fifo_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  fifo_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  fifo_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  fifo_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  fifo_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  fifo_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  fifo_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  fifo_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  fifo_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  fifo_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  fifo_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  fifo_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  fifo_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  fifo_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  fifo_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  fifo_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  fifo_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  fifo_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  fifo_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  fifo_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  fifo_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  fifo_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  fifo_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  fifo_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  fifo_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  fifo_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  fifo_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  fifo_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  fifo_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  fifo_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  fifo_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  fifo_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  fifo_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  fifo_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  fifo_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  fifo_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  fifo_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  fifo_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  fifo_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  fifo_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  fifo_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  fifo_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  fifo_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  fifo_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  fifo_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  fifo_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  fifo_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  fifo_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  fifo_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  fifo_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  fifo_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  fifo_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  fifo_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  fifo_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  fifo_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  fifo_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  fifo_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  fifo_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  fifo_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  fifo_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  fifo_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  fifo_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  fifo_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  fifo_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  fifo_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  fifo_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  fifo_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  fifo_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  fifo_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  fifo_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  fifo_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  fifo_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  fifo_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  fifo_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  fifo_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  fifo_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  fifo_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  fifo_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  fifo_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  fifo_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  fifo_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  fifo_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  fifo_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  fifo_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  fifo_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  fifo_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  fifo_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  fifo_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  fifo_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  fifo_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  fifo_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  fifo_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  fifo_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  fifo_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  fifo_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  fifo_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  fifo_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  fifo_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  fifo_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  fifo_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  fifo_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  fifo_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  fifo_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  fifo_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  fifo_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  fifo_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  fifo_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  fifo_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  fifo_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  fifo_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  fifo_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  fifo_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  fifo_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  fifo_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  fifo_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  fifo_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  fifo_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  fifo_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  fifo_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  fifo_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  fifo_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  fifo_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  fifo_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  fifo_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  fifo_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  fifo_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  fifo_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  fifo_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  fifo_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  fifo_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  fifo_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  fifo_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  fifo_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  fifo_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  fifo_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  fifo_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  fifo_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  fifo_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  fifo_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  fifo_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  fifo_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  fifo_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  fifo_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  fifo_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  fifo_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  fifo_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  fifo_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  fifo_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  fifo_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  fifo_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  fifo_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  fifo_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  fifo_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  fifo_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  fifo_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  fifo_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  fifo_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  fifo_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  fifo_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  fifo_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  fifo_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  fifo_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  fifo_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  fifo_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  fifo_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  fifo_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  fifo_255 = _RAND_255[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
